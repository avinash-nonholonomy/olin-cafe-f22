`timescale 1ns/1ps
`default_nettype none

module practice(rst, clk, ena, seed, out);

endmodule
