`timescale 1ns/1ps
`default_nettype none

module mux(in0, in1, select, out);

input in0, in1, select;
output logic out;

endmodule